-------------------------------------------------------------------------
-- Curt Lengemann
-------------------------------------------------------------------------


-- .vhd
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

package reg_package is
   
	type reg_array is array (31 downto 0) of std_logic_vector(31 downto 0);

end package reg_package;
 
-- Package Body Section
package body reg_package is

end package body reg_package;