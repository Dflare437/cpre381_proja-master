-------------------------------------------------------------------------
-- Curt Lengemann
-------------------------------------------------------------------------


-- tb_NBitALU.vhd
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_NBitALU is
    generic(N : integer := 32);
end tb_NBitALU;
    
architecture behavior of tb_NBitALU is


component NBit_ALU
    port(i_A : in std_logic_vector(N-1 downto 0);
	 i_B: in std_logic_vector(N-1 downto 0);
	 s_OPMUX : in std_logic_vector(3 downto 0);
	 ALU_Output: out std_logic_vector(N-1 downto 0);
	 o_ALUOverflow: out std_logic;
	 o_ALUCout: out std_logic;
	 o_ALUZero : out std_logic);
end component;

signal s_A, s_B, s_ALU_Output : std_logic_vector(N-1 downto 0);
signal signal_OPMUX : std_logic_vector(3 downto 0);
signal s_ALUOverflow, s_ALUCout, s_ALUZero : std_logic;

begin

DUT : NBit_ALU
	port map(i_A => s_A,
		 i_B => s_B,
		 s_OPMUX => signal_OPMUX,
		 ALU_Output => s_ALU_Output,
		 o_ALUOverflow => s_ALUOverflow,
		 o_ALUCout => s_ALUCout,
		 o_ALUZero => s_ALUZero);

P_TB: process
    begin

	--testing AND
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0000";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"00000000";
	signal_OPMUX <= "0000";
	wait for 100 ns;

	s_A <= x"00000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0000";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0000";
	wait for 100 ns;

	--testing OR
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0001";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"00000000";
	signal_OPMUX <= "0001";
	wait for 100 ns;

	s_A <= x"00000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0001";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0001";
	wait for 100 ns;

	--testing NOR
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0010";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"00000000";
	signal_OPMUX <= "0010";
	wait for 100 ns;

	s_A <= x"00000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0010";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0010";
	wait for 100 ns;

	--testing NAND
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0011";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"00000000";
	signal_OPMUX <= "0011";
	wait for 100 ns;

	s_A <= x"00000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0011";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0011";
	wait for 100 ns;

	--testing XOR
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0100";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"00000000";
	signal_OPMUX <= "0100";
	wait for 100 ns;

	s_A <= x"00000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0100";
	wait for 100 ns;

	s_A <= x"FFFFFFFF";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0100";
	wait for 100 ns;

	--testing ADD signed
	-- 2 positives
	s_A <= x"00000003";
	s_B <= x"00000006";
	signal_OPMUX <= "0101";
	wait for 100 ns;

	-- 2 negatives
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "0101";
	wait for 100 ns;

	-- one of each
	s_A <= x"0000000A";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "0101";
	wait for 100 ns;

	s_A <= x"FFFFFFFE";
	s_B <= x"0000000A";
	signal_OPMUX <= "0101";
	wait for 100 ns;

	--testing ADD unsigned
	-- 2 positives
	s_A <= x"00000003";
	s_B <= x"00000006";
	signal_OPMUX <= "1101";
	wait for 100 ns;

	-- 2 negatives
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "1101";
	wait for 100 ns;

	-- one of each
	s_A <= x"0000000A";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "1101";
	wait for 100 ns;

	s_A <= x"FFFFFFFE";
	s_B <= x"0000000A";
	signal_OPMUX <= "1101";
	wait for 100 ns;

	--testing SUB signed
	-- 2 positives
	s_A <= x"00000003";
	s_B <= x"00000006";
	signal_OPMUX <= "0110";
	wait for 100 ns;

	-- 2 negatives
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "0110";
	wait for 100 ns;

	-- one of each
	s_A <= x"0000000A";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "0110";
	wait for 100 ns;

	s_A <= x"FFFFFFFE";
	s_B <= x"0000000A";
	signal_OPMUX <= "0110";
	wait for 100 ns;

	--testing SUB unsigned
	-- 2 positives
	s_A <= x"00000003";
	s_B <= x"00000006";
	signal_OPMUX <= "1110";
	wait for 100 ns;

	-- 2 negatives
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "1110";
	wait for 100 ns;

	-- one of each
	s_A <= x"0000000A";
	s_B <= x"FFFFFFF9";
	signal_OPMUX <= "1110";
	wait for 100 ns;

	s_A <= x"FFFFFFFE";
	s_B <= x"0000000A";
	signal_OPMUX <= "1110";
	wait for 100 ns;

	-- testing SLT signed
	-- both positive LT
	s_A <= x"00000003";
	s_B <= x"00000009";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- both positive GT
	s_A <= x"00000009";
	s_B <= x"00000003";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- both negative LT
	s_A <= x"FFFFFFFD";
	s_B <= x"FFFFFFFE";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- both negative GT
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFFA";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- one of each LT
	s_A <= x"FFFFFFFB";
	s_B <= x"0000000C";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- one of each GT
	s_A <= x"00000003";
	s_B <= x"FFFFFFFE";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- both equal postive
	s_A <= x"00000003";
	s_B <= x"00000003";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- both equal negative
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFFE";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	--both 0
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	-- testing SLT unsigned
	-- both positive LT
	s_A <= x"00000003";
	s_B <= x"00000009";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- both positive GT
	s_A <= x"00000009";
	s_B <= x"00000003";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- both negative LT
	s_A <= x"FFFFFFFD";
	s_B <= x"FFFFFFFE";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- both negative GT
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFFA";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- one of each LT
	s_A <= x"FFFFFFFB";
	s_B <= x"0000000C";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- one of each GT
	s_A <= x"00000003";
	s_B <= x"FFFFFFFE";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- both equal postive
	s_A <= x"00000003";
	s_B <= x"00000003";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- both equal negative
	s_A <= x"FFFFFFFE";
	s_B <= x"FFFFFFFE";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	--both 0
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	--Testing edge cases
	--Overflow SLT signed
	s_A <= x"80000000";
	s_B <= x"7FFFFFFF";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	s_A <= x"7FFFFFFF";
	s_B <= x"80000000";
	signal_OPMUX <= "0111";
	wait for 100 ns;

	--Overflow SLT unsigned
	s_A <= x"80000000";
	s_B <= x"7FFFFFFF";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	s_A <= x"7FFFFFFF";
	s_B <= x"80000000";
	signal_OPMUX <= "1111";
	wait for 100 ns;

	-- Overflow add signed
	s_A <= x"00000001";
	s_B <= x"7FFFFFFF";
	signal_OPMUX <= "0101";
	wait for 100 ns;

	s_A <= x"80000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "0101";
	wait for 100 ns;

	-- Overflow add unsigned
	s_A <= x"00000001";
	s_B <= x"7FFFFFFF";
	signal_OPMUX <= "1101";
	wait for 100 ns;

	s_A <= x"80000000";
	s_B <= x"FFFFFFFF";
	signal_OPMUX <= "1101";
	wait for 100 ns;

	-- Overflow sub signed
	s_A <= x"FFFFFFFE";
	s_B <= x"7FFFFFFF";
	signal_OPMUX <= "0110";
	wait for 100 ns;

	s_A <= x"80000000";
	s_B <= x"00000001";
	signal_OPMUX <= "0110";
	wait for 100 ns;

	-- Overflow sub unsigned
	s_A <= x"FFFFFFFE";
	s_B <= x"7FFFFFFF";
	signal_OPMUX <= "1110";
	wait for 100 ns;

	s_A <= x"80000000";
	s_B <= x"00000001";
	signal_OPMUX <= "1110";
	wait for 100 ns;

	-- Check 0
	s_A <= x"00000000";
	s_B <= x"00000000";
	signal_OPMUX <= "0101";
	wait for 100 ns;


end process;
end behavior;